module gcd_fsm (
    input  logic clk,
    input logic rst,
    input logic go,
    input logic x_ne_y,
    input logic x_lt_y,
    output logic x_sel,
    output logic x_en,
    output logic y_sel,
    output logic y_en,
    output logic output_en,
    output logic done
);
  

// Your code here

endmodule